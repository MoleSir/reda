VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 2000 ;
END UNITS

MANUFACTURINGGRID 0.0050 ;

LAYER active
  TYPE MASTERSLICE ;
  MASK 1 ;
END active

LAYER nwell
  TYPE MASTERSLICE ;
  MASK 2 ;
END nwell

LAYER pwell
  TYPE MASTERSLICE ;
  MASK 3 ;
END pwell

LAYER nimplant
  TYPE MASTERSLICE ;
  MASK 4 ;
END nimplant

LAYER pimplant
  TYPE MASTERSLICE ;
  MASK 5 ;
END pimplant

LAYER poly
  TYPE MASTERSLICE ;
  MASK 9 ;
END poly

LAYER metal1
  TYPE ROUTING ;
  MASK 11 ;
  DIRECTION HORIZONTAL ;
  PITCH 0.13 ;
  WIDTH 0.065 ;
  AREA 0.0 ;
  SPACING 0.065 ;
END metal1

LAYER via1
  TYPE CUT ;
  MASK 12 ;
  SPACING 0.075 ;
  WIDTH 0.065 ;
  ENCLOSURE BELOW 0.035 0.035 ;
  ENCLOSURE ABOVE 0.035 0.035 ;
END via1

LAYER metal2
  TYPE ROUTING ;
  MASK 13 ;
  DIRECTION VERTICAL ;
  PITCH 0.14 ;
  WIDTH 0.07 ;
  AREA 0.0 ;
  SPACING 0.07 ;
END metal2

LAYER via2
  TYPE CUT ;
  MASK 14 ;
  SPACING 0.075 ;
  WIDTH 0.075 ;
  ENCLOSURE BELOW 0.035 0.035 ;
  ENCLOSURE ABOVE 0.035 0.035 ;
END via2

LAYER metal3
  TYPE ROUTING ;
  MASK 15 ;
  DIRECTION HORIZONTAL ;
  PITCH 0.14 ;
  WIDTH 0.07 ;
  AREA 0 ;
  SPACING 0.07 ;
END metal3

LAYER via3
  TYPE CUT ;
  MASK 16 ;
  SPACING 0.07 ;
  WIDTH 0.07 ;
  ENCLOSURE BELOW 0.035 0.035 ;
  ENCLOSURE ABOVE 0.035 0.035 ;
END via3

LAYER metal4
  TYPE ROUTING ;
  MASK 17 ;
  DIRECTION VERTICAL ;
  PITCH 0.14 ;
  WIDTH 0.14 ;
  AREA 0 ;
  SPACING 0.14 ;
END metal4

LAYER via4
  TYPE CUT ;
  MASK 18 ;
  SPACING 0.16 ;
  WIDTH 0.16 ;
  ENCLOSURE BELOW 0.03 0.03 ;
  ENCLOSURE ABOVE 0.03 0.03 ;
END via4

LAYER metal5
  TYPE ROUTING ;
  MASK 19 ;
  DIRECTION HORIZONTAL ;
  PITCH 0.14 ;
  WIDTH 0.14 ;
  AREA 0 ;
  SPACING 0.14 ;
END metal5

LAYER via5
  TYPE CUT ;
  MASK 20 ;
  SPACING 0.16 ;
  WIDTH 0.16 ;
  ENCLOSURE BELOW 0.03 0.03 ;
  ENCLOSURE ABOVE 0.03 0.03 ;
END via5

LAYER metal6
  TYPE ROUTING ;
  MASK 21 ;
  DIRECTION VERTICAL ;
  PITCH 0.14 ;
  WIDTH 0.14 ;
  AREA 0.017 ;
  SPACING 0.14 ;
END metal6

END LIBRARY
#
# End of file
#
